module drawGuess(clock, en, , counter, readPos, img, out);
  
endmodule